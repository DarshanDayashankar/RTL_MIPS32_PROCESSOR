`include "defines.v"

module ID_PIPE_EXE (CLK, RESET, DESTINATION_IN, REGISTER2_IN, OPERAND1_IN, OPERAND2_IN, PC_IN, OPERATOR_IN, 
                   MEM_READ_EN_IN, MEM_WRITE_EN_IN, WB_EN_IN, BRANCH_TAKEN_IN, SOURCE1_IN, SOURCE2_IN,
                   DESTINATION_OUT_REG, SW_OPERAND_OUT_REG, OPERAND1_OUT_REG, OPERAND2_OUT_REG, PC_OUT_REG,
                   OPERATOR_OUT_REG, MEM_READ_EN_OUT_REG, MEM_WRITE_EN_OUT_REG, WB_EN_OUT_REG, BRANCH_TAKEN_OUT_REG,
                   SOURCE1_OUT_REG, SOURCE2_OUT_REG);

    input CLK, RESET;
    input MEM_READ_EN_IN, MEM_WRITE_EN_IN, WB_EN_IN, BRANCH_TAKEN_IN;
    input [`OPERATOR_LEN-1:0] OPERATOR_IN;
    input [`WORD_LEN-1:0] REGISTER2_IN, OPERAND1_IN, OPERAND2_IN, PC_IN;
    input [`REG_ADDR_LEN-1:0] DESTINATION_IN, SOURCE1_IN, SOURCE2_IN;

    output reg MEM_READ_EN_OUT_REG, MEM_WRITE_EN_OUT_REG, WB_EN_OUT_REG, BRANCH_TAKEN_OUT_REG;
    output reg [`OPERATOR_LEN-1:0] OPERATOR_OUT_REG;
    output reg [`REG_ADDR_LEN-1:0] DESTINATION_OUT_REG, SOURCE1_OUT_REG, SOURCE2_OUT_REG;
    output reg [`WORD_LEN-1:0] SW_OPERAND_OUT_REG, OPERAND1_OUT_REG, OPERAND2_OUT_REG, PC_OUT_REG;

    always @ (posedge CLK) begin 
        if (RESET) begin 
            {MEM_READ_EN_OUT_REG, MEM_WRITE_EN_OUT_REG, WB_EN_OUT_REG, OPERATOR_OUT_REG, DESTINATION_OUT_REG, DESTINATION_OUT_REG,
            SW_OPERAND_OUT_REG, OPERAND1_OUT_REG, OPERAND2_OUT_REG, PC_OUT_REG, BRANCH_TAKEN_OUT_REG, SOURCE1_OUT_REG, SOURCE2_OUT_REG
            } <= 0;
        end
        else begin 
            MEM_READ_EN_OUT_REG <= MEM_READ_EN_IN;
            MEM_WRITE_EN_OUT_REG <= MEM_WRITE_EN_IN;
            WB_EN_OUT_REG <= MEM_READ_EN_IN;
            WB_EN_OUT_REG <= WB_EN_IN;
            OPERATOR_OUT_REG <= OPERATOR_IN;
            DESTINATION_OUT_REG <= DESTINATION_IN;
            SW_OPERAND_OUT_REG <= REGISTER2_IN;
            OPERAND1_OUT_REG <= OPERAND1_IN;
            OPERAND2_OUT_REG <= OPERAND2_IN;
            PC_OUT_REG <= PC_IN;
            BRANCH_TAKEN_OUT_REG <= BRANCH_TAKEN_IN;
            SOURCE1_OUT_REG <= SOURCE1_IN;
            SOURCE2_OUT_REG <= SOURCE2_IN; 
        end
    end

endmodule
