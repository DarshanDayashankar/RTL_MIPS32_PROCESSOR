`include "defines.v"

module INSTRUCTION_MEMORY (RESET, ADDRESS, INSTRUCTION);

parameter MEM_SIZE=`INSTR_MEM_SIZE;
input RESET;
input [`WORD_LEN-1:0] ADDRESS;
output reg [`WORD_LEN-1:0] INSTRUCTION;

wire [9:0] address = ADDRESS[9:0]; 

reg [`MEM_CELL_SIZE-1:0] MEM [0:MEM_SIZE-1];

always @ (ADDRESS) begin
    if (RESET == 1) begin
    
        MEM[0] <= 8'b10000000; //-- Addi	r1,r0,10
        MEM[1] <= 8'b00100000;
        MEM[2] <= 8'b00000000;
        MEM[3] <= 8'b00001010;

        MEM[4] <= 8'b00000100; //-- Add 	r2,r0,r1
        MEM[5] <= 8'b01000000;
        MEM[6] <= 8'b00001000;
        MEM[7] <= 8'b00000000;

        // MEM[8] <= 8'b00001100; //-- sub	r3,r0,r1
        // MEM[9] <= 8'b01100000;
        // MEM[10] <= 8'b00001000;
        // MEM[11] <= 8'b00000000;

        // MEM[12] <= 8'b00010100; //-- And	r4,r2,r3
        // MEM[13] <= 8'b10000010;
        // MEM[14] <= 8'b00011000;
        // MEM[15] <= 8'b00000000;

        // MEM[16] <= 8'b10000100; //-- Subi	r5,r0,564
        // MEM[17] <= 8'b10100000;
        // MEM[18] <= 8'b00000010;
        // MEM[19] <= 8'b00110100;

        // MEM[20] <= 8'b00011000; //-- or	r5,r5,r3
        // MEM[21] <= 8'b10100101;
        // MEM[22] <= 8'b00011000;
        // MEM[23] <= 8'b00000000;

        // MEM[24] <= 8'b00011100; //-- nor 	r6,r5,r0
        // MEM[25] <= 8'b11000101;
        // MEM[26] <= 8'b00000000;
        // MEM[27] <= 8'b00000000;

        // MEM[28] <= 8'b00100000; //-- xor	r0,r5,r1
        // MEM[29] <= 8'b00000101;
        // MEM[30] <= 8'b00001000;
        // MEM[31] <= 8'b00000000;

        // MEM[32] <= 8'b00100000; //-- xor	r7,r5,r0
        // MEM[33] <= 8'b11100101;
        // MEM[34] <= 8'b00001000;
        // MEM[35] <= 8'b00000000;

        // MEM[36] <= 8'b00100100; //-- sla	r7,r4,r2
        // MEM[37] <= 8'b11100100;
        // MEM[38] <= 8'b00010000;
        // MEM[39] <= 8'b00000000;

        // MEM[40] <= 8'b00101001; //-- sll	r8,r3,r2
        // MEM[41] <= 8'b00000011;
        // MEM[42] <= 8'b00010000;
        // MEM[43] <= 8'b00000000;

        // MEM[44] <= 8'b00101101; //-- sra	r9,r6,r2
        // MEM[45] <= 8'b00100110;
        // MEM[46] <= 8'b00010000;
        // MEM[47] <= 8'b00000000;

        // MEM[48] <= 8'b00110001; //-- srl	r10,r6,r2
        // MEM[49] <= 8'b01000110;
        // MEM[50] <= 8'b00010000;
        // MEM[51] <= 8'b00000000;

        // MEM[52] <= 8'b10000000; //-- Addi 	r1,r0,1024
        // MEM[53] <= 8'b00100000;
        // MEM[54] <= 8'b00000100;
        // MEM[55] <= 8'b00000000;

        // MEM[56] <= 8'b10010100; //-- st	r2,r1,0
        // MEM[57] <= 8'b01000001;
        // MEM[58] <= 8'b00000000;
        // MEM[59] <= 8'b00000000;

        // MEM[60] <= 8'b10010001; //-- ld	r11,r1,0
        // MEM[61] <= 8'b01100001;
        // MEM[62] <= 8'b00000000;
        // MEM[63] <= 8'b00000000;

        // MEM[64] <= 8'b10010100; //-- st	r3,r1,4
        // MEM[65] <= 8'b01100001;
        // MEM[66] <= 8'b00000000;
        // MEM[67] <= 8'b00000100;

        // MEM[68] <= 8'b10010100; //-- st	r4,r1,8
        // MEM[69] <= 8'b10000001;
        // MEM[70] <= 8'b00000000;
        // MEM[71] <= 8'b00001000;

        // MEM[72] <= 8'b10010100; //-- st	r5,r1,12
        // MEM[73] <= 8'b10100001;
        // MEM[74] <= 8'b00000000;
        // MEM[75] <= 8'b00001100;

        // MEM[76] <= 8'b10010100; //-- st	r6,r1,16
        // MEM[77] <= 8'b11000001;
        // MEM[78] <= 8'b00000000;
        // MEM[79] <= 8'b00010000;

        // MEM[80] <= 8'b10010100; //-- st	r7,r1,20
        // MEM[81] <= 8'b11100001;
        // MEM[82] <= 8'b00000000;
        // MEM[83] <= 8'b00010100;

        // MEM[84] <= 8'b10010101; //-- st	r8,r1,24
        // MEM[85] <= 8'b00000001;
        // MEM[86] <= 8'b00000000;
        // MEM[87] <= 8'b00011000;

        // MEM[88] <= 8'b10010101; //-- st	r9,r1,28
        // MEM[89] <= 8'b00100001;
        // MEM[90] <= 8'b00000000;
        // MEM[91] <= 8'b00011100;

        // MEM[92] <= 8'b10010101; //-- st	r10,r1,32
        // MEM[93] <= 8'b01000001;
        // MEM[94] <= 8'b00000000;
        // MEM[95] <= 8'b00100000;

        // MEM[96] <= 8'b10010101; //-- st	r11,r1,36
        // MEM[97] <= 8'b01100001;
        // MEM[98] <= 8'b00000000;
        // MEM[99] <= 8'b00100100;

        // MEM[100] <= 8'b10000000; //-- Addi 	r1,r0,3
        // MEM[101] <= 8'b00100000;
        // MEM[102] <= 8'b00000000;
        // MEM[103] <= 8'b00000011;

        // MEM[104] <= 8'b10000000; //-- Addi	r4,r0,1024
        // MEM[105] <= 8'b10000000;
        // MEM[106] <= 8'b00000100;
        // MEM[107] <= 8'b00000000;

        // MEM[108] <= 8'b10000000; //-- Addi 	r2,r0,0
        // MEM[109] <= 8'b01000000;
        // MEM[110] <= 8'b00000000;
        // MEM[111] <= 8'b00000000;

        // MEM[112] <= 8'b10000000; //-- Addi 	r3,r0,1
        // MEM[113] <= 8'b01100000;
        // MEM[114] <= 8'b00000000;
        // MEM[115] <= 8'b00000001;

        // MEM[116] <= 8'b10000001; //-- Addi 	r9,r0,2
        // MEM[117] <= 8'b00100000;
        // MEM[118] <= 8'b00000000;
        // MEM[119] <= 8'b00000010;

        // MEM[120] <= 8'b00101001; //-- sll	r8,r3,r9
        // MEM[121] <= 8'b00000011;
        // MEM[122] <= 8'b01001000;
        // MEM[123] <= 8'b00000000;

        // MEM[124] <= 8'b00000101; //-- Add 	r8,r4,r8
        // MEM[125] <= 8'b00000100;
        // MEM[126] <= 8'b01000000;
        // MEM[127] <= 8'b00000000;

        // MEM[128] <= 8'b10010000; //-- ld	r5,r8,0
        // MEM[129] <= 8'b10101000;
        // MEM[130] <= 8'b00000000;
        // MEM[131] <= 8'b00000000;

        // MEM[132] <= 8'b10010000; //-- ld	r6,r8,-4
        // MEM[133] <= 8'b11001000;
        // MEM[134] <= 8'b11111111;
        // MEM[135] <= 8'b11111100;

        // MEM[136] <= 8'b00001101; //-- sub 	r9,r5,r6
        // MEM[137] <= 8'b00100101;
        // MEM[138] <= 8'b00110000;
        // MEM[139] <= 8'b00000000;

        // MEM[140] <= 8'b10000001; //-- Addi 	r10,r0,0x8000
        // MEM[141] <= 8'b01000000;
        // MEM[142] <= 8'b10000000;
        // MEM[143] <= 8'b00000000;

        // MEM[144] <= 8'b10000001; //-- Addi	r11,r0,16
        // MEM[145] <= 8'b01100000;
        // MEM[146] <= 8'b00000000;
        // MEM[147] <= 8'b00010000;

        // MEM[148] <= 8'b00101001; //-- sll	r10,r10,r11
        // MEM[149] <= 8'b01001010;
        // MEM[150] <= 8'b01011000;
        // MEM[151] <= 8'b00000000;

        // MEM[152] <= 8'b00010101; //-- And 	r9,r9,r10
        // MEM[153] <= 8'b00101001;
        // MEM[154] <= 8'b01010000;
        // MEM[155] <= 8'b00000000;

        // MEM[156] <= 8'b10100000; //-- Bez	r9,2
        // MEM[157] <= 8'b00001001;
        // MEM[158] <= 8'b00000000;
        // MEM[159] <= 8'b00000010;

        // MEM[160] <= 8'b10010100; //-- st	r5,r8,-4
        // MEM[161] <= 8'b10101000;
        // MEM[162] <= 8'b11111111;
        // MEM[163] <= 8'b11111100;

        // MEM[164] <= 8'b10010100; //-- st	r6,r8,0
        // MEM[165] <= 8'b11001000;
        // MEM[166] <= 8'b00000000;
        // MEM[167] <= 8'b00000000;

        // MEM[168] <= 8'b10000000; //-- Addi 	r3,r3,1
        // MEM[169] <= 8'b01100011;
        // MEM[170] <= 8'b00000000;
        // MEM[171] <= 8'b00000001;

        // MEM[172] <= 8'b10100100; //-- BNE	r3,r1,-15
        // MEM[173] <= 8'b01100001;
        // MEM[174] <= 8'b11111111;
        // MEM[175] <= 8'b11110001;

        // MEM[176] <= 8'b10000000; //-- Addi 	r2,r2,1
        // MEM[177] <= 8'b01000010;
        // MEM[178] <= 8'b00000000;
        // MEM[179] <= 8'b00000001;

        // MEM[180] <= 8'b10100100; //-- BNE	r2,r1,-18
        // MEM[181] <= 8'b01000001;
        // MEM[182] <= 8'b11111111;
        // MEM[183] <= 8'b11101110;

        // MEM[184] <= 8'b10000000; //-- Addi 	r1,r0,1024
        // MEM[185] <= 8'b00100000;
        // MEM[186] <= 8'b00000100;
        // MEM[187] <= 8'b00000000;

        // MEM[188] <= 8'b10010000; //-- ld	r2,r1,0
        // MEM[189] <= 8'b01000001;
        // MEM[190] <= 8'b00000000;
        // MEM[191] <= 8'b00000000;

        // MEM[192] <= 8'b10010000; //-- ld	r3,r1,4
        // MEM[193] <= 8'b01100001;
        // MEM[194] <= 8'b00000000;
        // MEM[195] <= 8'b00000100;

        // MEM[196] <= 8'b10010000; //-- ld	r4,r1,8
        // MEM[197] <= 8'b10000001;
        // MEM[198] <= 8'b00000000;
        // MEM[199] <= 8'b00001000;

        // MEM[200] <= 8'b10010000; //-- ld	r5,r1,12
        // MEM[201] <= 8'b10100001;
        // MEM[202] <= 8'b00000000;
        // MEM[203] <= 8'b00001100;

        // MEM[204] <= 8'b10010000; //-- ld	r6,r1,16
        // MEM[205] <= 8'b11000001;
        // MEM[206] <= 8'b00000000;
        // MEM[207] <= 8'b00010000;

        // MEM[208] <= 8'b10010000; //-- ld	r7,r1,20
        // MEM[209] <= 8'b11100001;
        // MEM[210] <= 8'b00000000;
        // MEM[211] <= 8'b00010100;

        // MEM[212] <= 8'b10010001; //-- ld	r8,r1,24
        // MEM[213] <= 8'b00000001;
        // MEM[214] <= 8'b00000000;
        // MEM[215] <= 8'b00011000;

        // MEM[216] <= 8'b10010001; //-- ld	r9,r1,28
        // MEM[217] <= 8'b00100001;
        // MEM[218] <= 8'b00000000;
        // MEM[219] <= 8'b00011100;

        // MEM[220] <= 8'b10010001; //-- ld	r10,r1,32
        // MEM[221] <= 8'b01000001;
        // MEM[222] <= 8'b00000000;
        // MEM[223] <= 8'b00100000;

        // MEM[224] <= 8'b10010001; //-- ld	r11,r1,36
        // MEM[225] <= 8'b01100001;
        // MEM[226] <= 8'b00000000;
        // MEM[227] <= 8'b00100100;

        // MEM[228] <= 8'b10101000; //-- JMP 	-1
        // MEM[229] <= 8'b00000000;
        // MEM[230] <= 8'b11111111;
        // MEM[231] <= 8'b11111111;

        // MEM[232] <= 8'b00000000; //-- NOPE
        // MEM[233] <= 8'b00000000;
        // MEM[234] <= 8'b00000000;
        // MEM[235] <= 8'b00000000;
        
    end
    INSTRUCTION = {MEM[address], MEM[address + 1], MEM[address + 2], MEM[address + 3]};
end
endmodule 